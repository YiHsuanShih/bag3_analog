{{ _header }}

endmodule
